module top( in15 , in0 , in4 , in29 , in38 , in53 , in42 , in11 , in59 , in48 , in54 , in16 , in43 , in37 , in61 , in14 , in62 , in60 , in40 , in5 , in28 , in7 , in6 , in34 , in57 , in3 , in56 , in45 , in10 , in27 , in21 , in25 , in22 , in12 , in58 , in36 , in51 , in18 , in9 , in39 , in24 , in26 , in8 , in41 , in55 , in2 , in49 , in19 , in35 , in50 , in32 , in30 , in33 , in17 , in31 , in44 , in1 , in23 , in52 , in20 , in46 , in13 , in63 , in47 , out1 , out3 , out6 , out2 , out4 , out5 );
  input in15 , in0 , in4 , in29 , in38 , in53 , in42 , in11 , in59 , in48 , in54 , in16 , in43 , in37 , in61 , in14 , in62 , in60 , in40 , in5 , in28 , in7 , in6 , in34 , in57 , in3 , in56 , in45 , in10 , in27 , in21 , in25 , in22 , in12 , in58 , in36 , in51 , in18 , in9 , in39 , in24 , in26 , in8 , in41 , in55 , in2 , in49 , in19 , in35 , in50 , in32 , in30 , in33 , in17 , in31 , in44 , in1 , in23 , in52 , in20 , in46 , in13 , in63 , in47 ;
  output out1 , out3 , out6 , out2 , out4 , out5 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 ;
  assign n65 = in15 & in14 ;
  assign n66 = in12 | in13 ;
  assign n67 = in4 | in5 ;
  assign n68 = in0 | in1 ;
  assign n69 = in3 & in2 ;
  assign n70 = ( n67 & n68 ) | ( n67 & n69 ) | ( n68 & n69 ) ;
  assign n71 = ( ~n67 & n68 ) | ( ~n67 & n69 ) | ( n68 & n69 ) ;
  assign n72 = ( n67 & ~n70 ) | ( n67 & n71 ) | ( ~n70 & n71 ) ;
  assign n73 = in11 & in10 ;
  assign n74 = in7 & in6 ;
  assign n75 = in9 | in8 ;
  assign n76 = ( n73 & n74 ) | ( n73 & n75 ) | ( n74 & n75 ) ;
  assign n77 = ( ~n73 & n74 ) | ( ~n73 & n75 ) | ( n74 & n75 ) ;
  assign n78 = ( n73 & ~n76 ) | ( n73 & n77 ) | ( ~n76 & n77 ) ;
  assign n79 = ( n66 & n72 ) | ( n66 & n78 ) | ( n72 & n78 ) ;
  assign n80 = ( ~n66 & n72 ) | ( ~n66 & n78 ) | ( n72 & n78 ) ;
  assign n81 = ( n66 & ~n79 ) | ( n66 & n80 ) | ( ~n79 & n80 ) ;
  assign n82 = n65 & n81 ;
  assign n83 = n65 | n81 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = in30 & in31 ;
  assign n86 = in29 | in28 ;
  assign n87 = in21 | in20 ;
  assign n88 = in16 | in17 ;
  assign n89 = in18 & in19 ;
  assign n90 = ( n87 & n88 ) | ( n87 & n89 ) | ( n88 & n89 ) ;
  assign n91 = ( ~n87 & n88 ) | ( ~n87 & n89 ) | ( n88 & n89 ) ;
  assign n92 = ( n87 & ~n90 ) | ( n87 & n91 ) | ( ~n90 & n91 ) ;
  assign n93 = in27 & in26 ;
  assign n94 = in22 & in23 ;
  assign n95 = in25 | in24 ;
  assign n96 = ( n93 & n94 ) | ( n93 & n95 ) | ( n94 & n95 ) ;
  assign n97 = ( ~n93 & n94 ) | ( ~n93 & n95 ) | ( n94 & n95 ) ;
  assign n98 = ( n93 & ~n96 ) | ( n93 & n97 ) | ( ~n96 & n97 ) ;
  assign n99 = ( n86 & n92 ) | ( n86 & n98 ) | ( n92 & n98 ) ;
  assign n100 = ( ~n86 & n92 ) | ( ~n86 & n98 ) | ( n92 & n98 ) ;
  assign n101 = ( n86 & ~n99 ) | ( n86 & n100 ) | ( ~n99 & n100 ) ;
  assign n102 = n85 & n101 ;
  assign n103 = n85 | n101 ;
  assign n104 = ~n102 & n103 ;
  assign n105 = n84 & n104 ;
  assign n106 = n84 | n104 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = in46 & in47 ;
  assign n109 = in45 | in44 ;
  assign n110 = in37 | in36 ;
  assign n111 = in32 | in33 ;
  assign n112 = in34 & in35 ;
  assign n113 = ( n110 & n111 ) | ( n110 & n112 ) | ( n111 & n112 ) ;
  assign n114 = ( ~n110 & n111 ) | ( ~n110 & n112 ) | ( n111 & n112 ) ;
  assign n115 = ( n110 & ~n113 ) | ( n110 & n114 ) | ( ~n113 & n114 ) ;
  assign n116 = in42 & in43 ;
  assign n117 = in38 & in39 ;
  assign n118 = in40 | in41 ;
  assign n119 = ( n116 & n117 ) | ( n116 & n118 ) | ( n117 & n118 ) ;
  assign n120 = ( ~n116 & n117 ) | ( ~n116 & n118 ) | ( n117 & n118 ) ;
  assign n121 = ( n116 & ~n119 ) | ( n116 & n120 ) | ( ~n119 & n120 ) ;
  assign n122 = ( n109 & n115 ) | ( n109 & n121 ) | ( n115 & n121 ) ;
  assign n123 = ( ~n109 & n115 ) | ( ~n109 & n121 ) | ( n115 & n121 ) ;
  assign n124 = ( n109 & ~n122 ) | ( n109 & n123 ) | ( ~n122 & n123 ) ;
  assign n125 = n108 & n124 ;
  assign n126 = n108 | n124 ;
  assign n127 = ~n125 & n126 ;
  assign n128 = in62 & in63 ;
  assign n129 = in61 | in60 ;
  assign n130 = in53 | in52 ;
  assign n131 = in48 | in49 ;
  assign n132 = in51 & in50 ;
  assign n133 = ( n130 & n131 ) | ( n130 & n132 ) | ( n131 & n132 ) ;
  assign n134 = ( ~n130 & n131 ) | ( ~n130 & n132 ) | ( n131 & n132 ) ;
  assign n135 = ( n130 & ~n133 ) | ( n130 & n134 ) | ( ~n133 & n134 ) ;
  assign n136 = in59 & in58 ;
  assign n137 = in54 & in55 ;
  assign n138 = in57 | in56 ;
  assign n139 = ( n136 & n137 ) | ( n136 & n138 ) | ( n137 & n138 ) ;
  assign n140 = ( ~n136 & n137 ) | ( ~n136 & n138 ) | ( n137 & n138 ) ;
  assign n141 = ( n136 & ~n139 ) | ( n136 & n140 ) | ( ~n139 & n140 ) ;
  assign n142 = ( n129 & n135 ) | ( n129 & n141 ) | ( n135 & n141 ) ;
  assign n143 = ( ~n129 & n135 ) | ( ~n129 & n141 ) | ( n135 & n141 ) ;
  assign n144 = ( n129 & ~n142 ) | ( n129 & n143 ) | ( ~n142 & n143 ) ;
  assign n145 = n128 | n144 ;
  assign n146 = n128 & n144 ;
  assign n147 = n145 & ~n146 ;
  assign n148 = n127 & n147 ;
  assign n149 = n127 | n147 ;
  assign n150 = ~n148 & n149 ;
  assign n151 = n107 & n150 ;
  assign n152 = n107 | n150 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = ( n70 & n76 ) | ( n70 & n79 ) | ( n76 & n79 ) ;
  assign n155 = ( n70 & n76 ) | ( n70 & ~n79 ) | ( n76 & ~n79 ) ;
  assign n156 = ( n79 & ~n154 ) | ( n79 & n155 ) | ( ~n154 & n155 ) ;
  assign n157 = n82 & n156 ;
  assign n158 = n154 & n157 ;
  assign n159 = n154 | n157 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = ( n90 & n96 ) | ( n90 & n99 ) | ( n96 & n99 ) ;
  assign n162 = ( n90 & n96 ) | ( n90 & ~n99 ) | ( n96 & ~n99 ) ;
  assign n163 = ( n99 & ~n161 ) | ( n99 & n162 ) | ( ~n161 & n162 ) ;
  assign n164 = n102 & n163 ;
  assign n165 = n161 & n164 ;
  assign n166 = n161 | n164 ;
  assign n167 = ~n165 & n166 ;
  assign n168 = n160 & n167 ;
  assign n169 = n160 | n167 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = n82 | n156 ;
  assign n172 = ~n157 & n171 ;
  assign n173 = n102 | n163 ;
  assign n174 = ~n164 & n173 ;
  assign n175 = ( n105 & n172 ) | ( n105 & n174 ) | ( n172 & n174 ) ;
  assign n176 = n170 & n175 ;
  assign n177 = n170 | n175 ;
  assign n178 = ~n176 & n177 ;
  assign n179 = ( n113 & n119 ) | ( n113 & n122 ) | ( n119 & n122 ) ;
  assign n180 = ( n113 & n119 ) | ( n113 & ~n122 ) | ( n119 & ~n122 ) ;
  assign n181 = ( n122 & ~n179 ) | ( n122 & n180 ) | ( ~n179 & n180 ) ;
  assign n182 = n125 & n181 ;
  assign n183 = n179 & n182 ;
  assign n184 = n179 | n182 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = ( n133 & n139 ) | ( n133 & n142 ) | ( n139 & n142 ) ;
  assign n187 = ( n133 & n139 ) | ( n133 & ~n142 ) | ( n139 & ~n142 ) ;
  assign n188 = ( n142 & ~n186 ) | ( n142 & n187 ) | ( ~n186 & n187 ) ;
  assign n189 = n146 & n188 ;
  assign n190 = n186 & n189 ;
  assign n191 = n186 | n189 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = n185 & n192 ;
  assign n194 = n185 | n192 ;
  assign n195 = ~n193 & n194 ;
  assign n196 = n125 | n181 ;
  assign n197 = ~n182 & n196 ;
  assign n198 = n146 | n188 ;
  assign n199 = ~n189 & n198 ;
  assign n200 = ( n148 & n197 ) | ( n148 & n199 ) | ( n197 & n199 ) ;
  assign n201 = n195 & n200 ;
  assign n202 = n195 | n200 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = n178 & n203 ;
  assign n205 = n178 | n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = n172 & n174 ;
  assign n208 = n172 | n174 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = n105 & n209 ;
  assign n211 = n105 | n209 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n197 & n199 ;
  assign n214 = n197 | n199 ;
  assign n215 = ~n213 & n214 ;
  assign n216 = n148 & n215 ;
  assign n217 = n148 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ( n151 & n212 ) | ( n151 & n218 ) | ( n212 & n218 ) ;
  assign n220 = n206 & n219 ;
  assign n221 = n206 | n219 ;
  assign n222 = ~n220 & n221 ;
  assign n223 = ( n160 & n167 ) | ( n160 & n175 ) | ( n167 & n175 ) ;
  assign n224 = ( n158 & n165 ) | ( n158 & n223 ) | ( n165 & n223 ) ;
  assign n225 = ( n185 & n192 ) | ( n185 & n200 ) | ( n192 & n200 ) ;
  assign n226 = ( n183 & n190 ) | ( n183 & n225 ) | ( n190 & n225 ) ;
  assign n227 = n158 & n165 ;
  assign n228 = n158 | n165 ;
  assign n229 = ~n227 & n228 ;
  assign n230 = n223 & n229 ;
  assign n231 = n223 | n229 ;
  assign n232 = ~n230 & n231 ;
  assign n233 = n183 & n190 ;
  assign n234 = n183 | n190 ;
  assign n235 = ~n233 & n234 ;
  assign n236 = n225 & n235 ;
  assign n237 = n225 | n235 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ( n178 & n203 ) | ( n178 & n219 ) | ( n203 & n219 ) ;
  assign n240 = ( n232 & n238 ) | ( n232 & n239 ) | ( n238 & n239 ) ;
  assign n241 = ( n224 & n226 ) | ( n224 & n240 ) | ( n226 & n240 ) ;
  assign n242 = n212 & n218 ;
  assign n243 = n212 | n218 ;
  assign n244 = ~n242 & n243 ;
  assign n245 = n151 & n244 ;
  assign n246 = n151 | n244 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = n232 & n238 ;
  assign n249 = n232 | n238 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = n239 & n250 ;
  assign n252 = n239 | n250 ;
  assign n253 = ~n251 & n252 ;
  assign n254 = n224 & n226 ;
  assign n255 = n224 | n226 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = n240 & n256 ;
  assign n258 = n240 | n256 ;
  assign n259 = ~n257 & n258 ;
  assign out1 = n153 ;
  assign out3 = n222 ;
  assign out6 = n241 ;
  assign out2 = n247 ;
  assign out4 = n253 ;
  assign out5 = n259 ;
endmodule
