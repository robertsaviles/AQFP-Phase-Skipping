module top( in0 , in1 , in2 , in3 , in4 , in5 , in6 , in7 , in8 , in9 , in10 , in11 , in12 , in13 , in14 , in15 , out1 , out2 , out3 , out4 );
  input in0 , in1 , in2 , in3 , in4 , in5 , in6 , in7 , in8 , in9 , in10 , in11 , in12 , in13 , in14 , in15 ;
  output out1 , out2 , out3 , out4 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n17 = in14 & in15 ;
  assign n18 = in12 | in13 ;
  assign n19 = in4 | in5 ;
  assign n20 = in0 | in1 ;
  assign n21 = in2 & in3 ;
  assign n22 = ( n19 & n20 ) | ( n19 & n21 ) | ( n20 & n21 ) ;
  assign n23 = ( ~n19 & n20 ) | ( ~n19 & n21 ) | ( n20 & n21 ) ;
  assign n24 = ( n19 & ~n22 ) | ( n19 & n23 ) | ( ~n22 & n23 ) ;
  assign n25 = in10 & in11 ;
  assign n26 = in6 & in7 ;
  assign n27 = in8 | in9 ;
  assign n28 = ( n25 & n26 ) | ( n25 & n27 ) | ( n26 & n27 ) ;
  assign n29 = ( ~n25 & n26 ) | ( ~n25 & n27 ) | ( n26 & n27 ) ;
  assign n30 = ( n25 & ~n28 ) | ( n25 & n29 ) | ( ~n28 & n29 ) ;
  assign n31 = ( n18 & n24 ) | ( n18 & n30 ) | ( n24 & n30 ) ;
  assign n32 = ( ~n18 & n24 ) | ( ~n18 & n30 ) | ( n24 & n30 ) ;
  assign n33 = ( n18 & ~n31 ) | ( n18 & n32 ) | ( ~n31 & n32 ) ;
  assign n34 = n17 & n33 ;
  assign n35 = n17 | n33 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = ( n22 & n28 ) | ( n22 & n31 ) | ( n28 & n31 ) ;
  assign n38 = ( n22 & n28 ) | ( n22 & ~n31 ) | ( n28 & ~n31 ) ;
  assign n39 = ( n31 & ~n37 ) | ( n31 & n38 ) | ( ~n37 & n38 ) ;
  assign n40 = n34 & n39 ;
  assign n41 = n34 | n39 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n37 & n40 ;
  assign n44 = n37 | n40 ;
  assign n45 = ~n43 & n44 ;
  assign out1 = n36 ;
  assign out2 = n42 ;
  assign out3 = n45 ;
  assign out4 = n43 ;
endmodule
