module top( in6 , in15 , in13 , in14 , in2 , in10 , in24 , in8 , in22 , in20 , in7 , in25 , in5 , in4 , in23 , in27 , in1 , in0 , in16 , in30 , in26 , in12 , in11 , in17 , in19 , in18 , in21 , in31 , in29 , in28 , in9 , in3 , out2 , out1 , out3 , out5 , out4 );
  input in6 , in15 , in13 , in14 , in2 , in10 , in24 , in8 , in22 , in20 , in7 , in25 , in5 , in4 , in23 , in27 , in1 , in0 , in16 , in30 , in26 , in12 , in11 , in17 , in19 , in18 , in21 , in31 , in29 , in28 , in9 , in3 ;
  output out2 , out1 , out3 , out5 , out4 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ;
  assign n33 = in29 | in28 ;
  assign n34 = in20 | in21 ;
  assign n35 = in16 | in17 ;
  assign n36 = in19 & in18 ;
  assign n37 = ( n34 & n35 ) | ( n34 & n36 ) | ( n35 & n36 ) ;
  assign n38 = ( ~n34 & n35 ) | ( ~n34 & n36 ) | ( n35 & n36 ) ;
  assign n39 = ( n34 & ~n37 ) | ( n34 & n38 ) | ( ~n37 & n38 ) ;
  assign n40 = in27 & in26 ;
  assign n41 = in22 & in23 ;
  assign n42 = in24 | in25 ;
  assign n43 = ( n40 & n41 ) | ( n40 & n42 ) | ( n41 & n42 ) ;
  assign n44 = ( ~n40 & n41 ) | ( ~n40 & n42 ) | ( n41 & n42 ) ;
  assign n45 = ( n40 & ~n43 ) | ( n40 & n44 ) | ( ~n43 & n44 ) ;
  assign n46 = ( n33 & n39 ) | ( n33 & n45 ) | ( n39 & n45 ) ;
  assign n47 = ( n37 & n43 ) | ( n37 & n46 ) | ( n43 & n46 ) ;
  assign n48 = ( n37 & n43 ) | ( n37 & ~n46 ) | ( n43 & ~n46 ) ;
  assign n49 = ( n46 & ~n47 ) | ( n46 & n48 ) | ( ~n47 & n48 ) ;
  assign n50 = in30 & in31 ;
  assign n51 = ( ~n33 & n39 ) | ( ~n33 & n45 ) | ( n39 & n45 ) ;
  assign n52 = ( n33 & ~n46 ) | ( n33 & n51 ) | ( ~n46 & n51 ) ;
  assign n53 = n50 & n52 ;
  assign n54 = n49 & n53 ;
  assign n55 = n49 | n53 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = in13 | in12 ;
  assign n58 = in5 | in4 ;
  assign n59 = in1 | in0 ;
  assign n60 = in2 & in3 ;
  assign n61 = ( n58 & n59 ) | ( n58 & n60 ) | ( n59 & n60 ) ;
  assign n62 = ( ~n58 & n59 ) | ( ~n58 & n60 ) | ( n59 & n60 ) ;
  assign n63 = ( n58 & ~n61 ) | ( n58 & n62 ) | ( ~n61 & n62 ) ;
  assign n64 = in10 & in11 ;
  assign n65 = in6 & in7 ;
  assign n66 = in8 | in9 ;
  assign n67 = ( n64 & n65 ) | ( n64 & n66 ) | ( n65 & n66 ) ;
  assign n68 = ( ~n64 & n65 ) | ( ~n64 & n66 ) | ( n65 & n66 ) ;
  assign n69 = ( n64 & ~n67 ) | ( n64 & n68 ) | ( ~n67 & n68 ) ;
  assign n70 = ( n57 & n63 ) | ( n57 & n69 ) | ( n63 & n69 ) ;
  assign n71 = ( n61 & n67 ) | ( n61 & n70 ) | ( n67 & n70 ) ;
  assign n72 = ( n61 & n67 ) | ( n61 & ~n70 ) | ( n67 & ~n70 ) ;
  assign n73 = ( n70 & ~n71 ) | ( n70 & n72 ) | ( ~n71 & n72 ) ;
  assign n74 = in15 & in14 ;
  assign n75 = ( ~n57 & n63 ) | ( ~n57 & n69 ) | ( n63 & n69 ) ;
  assign n76 = ( n57 & ~n70 ) | ( n57 & n75 ) | ( ~n70 & n75 ) ;
  assign n77 = n74 & n76 ;
  assign n78 = n73 & n77 ;
  assign n79 = n73 | n77 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = n56 & n80 ;
  assign n82 = n56 | n80 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = n50 | n52 ;
  assign n85 = ~n53 & n84 ;
  assign n86 = n74 | n76 ;
  assign n87 = ~n77 & n86 ;
  assign n88 = n85 & n87 ;
  assign n89 = n83 & n88 ;
  assign n90 = n83 | n88 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = n85 | n87 ;
  assign n93 = ~n88 & n92 ;
  assign n94 = n47 & n54 ;
  assign n95 = n47 | n54 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = n71 & n78 ;
  assign n98 = n71 | n78 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = n96 & n99 ;
  assign n101 = n96 | n99 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = ( n56 & n80 ) | ( n56 & n88 ) | ( n80 & n88 ) ;
  assign n104 = n102 & n103 ;
  assign n105 = n102 | n103 ;
  assign n106 = ~n104 & n105 ;
  assign n107 = ( n96 & n99 ) | ( n96 & n103 ) | ( n99 & n103 ) ;
  assign n108 = ( n94 & n97 ) | ( n94 & n107 ) | ( n97 & n107 ) ;
  assign n109 = n94 | n97 ;
  assign n110 = n94 & n97 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = n107 & n111 ;
  assign n113 = n107 | n111 ;
  assign n114 = ~n112 & n113 ;
  assign out2 = n91 ;
  assign out1 = n93 ;
  assign out3 = n106 ;
  assign out5 = n108 ;
  assign out4 = n114 ;
endmodule
