module top( ioin21 , ioin17 , ioin24 , ioin216 , ioin111 , ioin226 , iofn0 , ioin212 , ioin221 , ioin214 , ioin13 , ioin117 , ioin120 , ioin16 , ioin15 , ioin118 , ioin227 , ioin228 , ioin225 , ioin114 , ioin217 , ioin125 , ioin12 , ioin115 , ioin222 , ioin18 , ioin121 , ioin223 , ioin119 , ioin26 , ioin29 , ioin23 , ioin113 , ioin123 , ioin213 , ioin112 , ioin10 , ioin215 , iofn2 , ioin128 , ioin28 , ioin131 , ioin20 , ioin220 , ioin25 , ioin229 , ioin231 , ioin218 , ioin116 , ioin11 , ioin129 , ioin224 , ioin230 , ioin19 , ioin130 , ioin219 , ioin27 , ioin22 , ioin127 , ioin211 , ioin124 , iofn3 , ioin210 , iofn1 , ioin14 , ioin126 , ioin110 , ioin122 , ioout22 , ioadderout22 , ioout7 , iotestadderCout , ioadderout17 , ioadderout26 , ioadderout1 , ioadderout23 , ioout1 , ioadderout8 , ioadderout0 , ioadderout7 , ioout15 , ioout31 , ioadderout10 , ioout25 , ioout10 , ioout14 , ioout24 , ioadderout5 , ioout12 , ioadderout9 , ioadderout30 , ioadderout12 , ioadderout13 , ioout13 , ioout21 , ioadderout16 , ioout30 , ioadderout2 , ioout2 , ioadderout31 , ioadderout14 , ioout26 , ioout17 , ioadderout6 , ioout18 , ioout0 , ioout4 , ioout19 , ioadderout19 , ioout23 , ioout8 , ioadderout20 , ioout20 , ioadderout25 , ioadderout29 , ioadderout15 , ioout3 , ioout28 , ioout27 , ioadderout11 , ioout5 , ioadderout4 , ioout9 , ioadderout28 , ioadderout21 , ioadderout24 , ioout29 , ioadderout27 , ioout16 , ioout11 , ioout6 , ioadderout3 , ioadderout18 );
  input ioin21 , ioin17 , ioin24 , ioin216 , ioin111 , ioin226 , iofn0 , ioin212 , ioin221 , ioin214 , ioin13 , ioin117 , ioin120 , ioin16 , ioin15 , ioin118 , ioin227 , ioin228 , ioin225 , ioin114 , ioin217 , ioin125 , ioin12 , ioin115 , ioin222 , ioin18 , ioin121 , ioin223 , ioin119 , ioin26 , ioin29 , ioin23 , ioin113 , ioin123 , ioin213 , ioin112 , ioin10 , ioin215 , iofn2 , ioin128 , ioin28 , ioin131 , ioin20 , ioin220 , ioin25 , ioin229 , ioin231 , ioin218 , ioin116 , ioin11 , ioin129 , ioin224 , ioin230 , ioin19 , ioin130 , ioin219 , ioin27 , ioin22 , ioin127 , ioin211 , ioin124 , iofn3 , ioin210 , iofn1 , ioin14 , ioin126 , ioin110 , ioin122 ;
  output ioout22 , ioadderout22 , ioout7 , iotestadderCout , ioadderout17 , ioadderout26 , ioadderout1 , ioadderout23 , ioout1 , ioadderout8 , ioadderout0 , ioadderout7 , ioout15 , ioout31 , ioadderout10 , ioout25 , ioout10 , ioout14 , ioout24 , ioadderout5 , ioout12 , ioadderout9 , ioadderout30 , ioadderout12 , ioadderout13 , ioout13 , ioout21 , ioadderout16 , ioout30 , ioadderout2 , ioout2 , ioadderout31 , ioadderout14 , ioout26 , ioout17 , ioadderout6 , ioout18 , ioout0 , ioout4 , ioout19 , ioadderout19 , ioout23 , ioout8 , ioadderout20 , ioout20 , ioadderout25 , ioadderout29 , ioadderout15 , ioout3 , ioout28 , ioout27 , ioadderout11 , ioout5 , ioadderout4 , ioout9 , ioadderout28 , ioadderout21 , ioadderout24 , ioout29 , ioadderout27 , ioout16 , ioout11 , ioout6 , ioadderout3 , ioadderout18 ;
  wire n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 ;
  assign n69 = ~iofn0 & iofn3 ;
  assign n70 = ~iofn2 & iofn1 ;
  assign n71 = n69 & n70 ;
  assign n72 = iofn2 | iofn3 ;
  assign n73 = iofn0 | iofn1 ;
  assign n74 = n72 | n73 ;
  assign n75 = ~n71 & n74 ;
  assign n76 = ioin21 | ioin20 ;
  assign n77 = ioin22 | n76 ;
  assign n78 = ioin23 | n77 ;
  assign n79 = ioin24 | n78 ;
  assign n80 = ioin25 | n79 ;
  assign n81 = ioin26 | n80 ;
  assign n82 = ioin27 | n81 ;
  assign n83 = ioin28 | n82 ;
  assign n84 = ioin29 | n83 ;
  assign n85 = ioin210 | n84 ;
  assign n86 = ioin211 | n85 ;
  assign n87 = ioin212 | n86 ;
  assign n88 = ioin213 | n87 ;
  assign n89 = ioin214 | n88 ;
  assign n90 = ioin215 | n89 ;
  assign n91 = ioin216 | n90 ;
  assign n92 = ioin217 | n91 ;
  assign n93 = ioin218 | n92 ;
  assign n94 = ioin219 | n93 ;
  assign n95 = ioin220 | n94 ;
  assign n96 = ioin221 | n95 ;
  assign n97 = iofn3 & n96 ;
  assign n98 = ~ioin222 & n97 ;
  assign n99 = ioin222 & ~n97 ;
  assign n100 = n98 | n99 ;
  assign n101 = ioin10 & ioin20 ;
  assign n102 = ioin11 | n101 ;
  assign n103 = ioin11 & n101 ;
  assign n104 = ioin21 & ~iofn3 ;
  assign n105 = ioin21 & ioin20 ;
  assign n106 = iofn3 & n76 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = n104 | n107 ;
  assign n109 = n103 | n108 ;
  assign n110 = n102 & n109 ;
  assign n111 = ioin12 | n110 ;
  assign n112 = ioin12 & n110 ;
  assign n113 = ~ioin22 & n106 ;
  assign n114 = ioin22 & ~n106 ;
  assign n115 = n113 | n114 ;
  assign n116 = n112 | n115 ;
  assign n117 = n111 & n116 ;
  assign n118 = ioin13 | n117 ;
  assign n119 = ioin13 & n117 ;
  assign n120 = iofn3 & n77 ;
  assign n121 = ioin23 & n120 ;
  assign n122 = ioin23 | n120 ;
  assign n123 = ~n121 & n122 ;
  assign n124 = n119 | n123 ;
  assign n125 = n118 & n124 ;
  assign n126 = ioin14 | n125 ;
  assign n127 = ioin14 & n125 ;
  assign n128 = iofn3 & n78 ;
  assign n129 = ~ioin24 & n128 ;
  assign n130 = ioin24 & ~n128 ;
  assign n131 = n129 | n130 ;
  assign n132 = n127 | n131 ;
  assign n133 = n126 & n132 ;
  assign n134 = ioin15 | n133 ;
  assign n135 = ioin15 & n133 ;
  assign n136 = iofn3 & n79 ;
  assign n137 = ioin25 & n136 ;
  assign n138 = ioin25 | n136 ;
  assign n139 = ~n137 & n138 ;
  assign n140 = n135 | n139 ;
  assign n141 = n134 & n140 ;
  assign n142 = ioin16 & n141 ;
  assign n143 = ioin16 | n141 ;
  assign n144 = iofn3 & n80 ;
  assign n145 = ~ioin26 & n144 ;
  assign n146 = ioin26 & ~n144 ;
  assign n147 = n145 | n146 ;
  assign n148 = n143 & n147 ;
  assign n149 = n142 | n148 ;
  assign n150 = ioin17 | n149 ;
  assign n151 = ioin17 & n149 ;
  assign n152 = iofn3 & n81 ;
  assign n153 = ioin27 & n152 ;
  assign n154 = ioin27 | n152 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = n151 | n155 ;
  assign n157 = n150 & n156 ;
  assign n158 = ioin18 | n157 ;
  assign n159 = ioin18 & n157 ;
  assign n160 = iofn3 & n82 ;
  assign n161 = ~ioin28 & n160 ;
  assign n162 = ioin28 & ~n160 ;
  assign n163 = n161 | n162 ;
  assign n164 = n159 | n163 ;
  assign n165 = n158 & n164 ;
  assign n166 = ioin19 | n165 ;
  assign n167 = iofn3 & n83 ;
  assign n168 = ioin29 & n167 ;
  assign n169 = ioin29 | n167 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = ioin19 & n165 ;
  assign n172 = n170 | n171 ;
  assign n173 = n166 & n172 ;
  assign n174 = ioin110 | n173 ;
  assign n175 = iofn3 & n84 ;
  assign n176 = ~ioin210 & n175 ;
  assign n177 = ioin210 & ~n175 ;
  assign n178 = n176 | n177 ;
  assign n179 = ioin110 & n173 ;
  assign n180 = n178 | n179 ;
  assign n181 = n174 & n180 ;
  assign n182 = ioin111 | n181 ;
  assign n183 = iofn3 & n85 ;
  assign n184 = ioin211 & n183 ;
  assign n185 = ioin211 | n183 ;
  assign n186 = ~n184 & n185 ;
  assign n187 = ioin111 & n181 ;
  assign n188 = n186 | n187 ;
  assign n189 = n182 & n188 ;
  assign n190 = ioin112 | n189 ;
  assign n191 = iofn3 & n86 ;
  assign n192 = ~ioin212 & n191 ;
  assign n193 = ioin212 & ~n191 ;
  assign n194 = n192 | n193 ;
  assign n195 = ioin112 & n189 ;
  assign n196 = n194 | n195 ;
  assign n197 = n190 & n196 ;
  assign n198 = ioin113 | n197 ;
  assign n199 = iofn3 & n87 ;
  assign n200 = ioin213 & n199 ;
  assign n201 = ioin213 | n199 ;
  assign n202 = ~n200 & n201 ;
  assign n203 = ioin113 & n197 ;
  assign n204 = n202 | n203 ;
  assign n205 = n198 & n204 ;
  assign n206 = ioin114 | n205 ;
  assign n207 = iofn3 & n88 ;
  assign n208 = ~ioin214 & n207 ;
  assign n209 = ioin214 & ~n207 ;
  assign n210 = n208 | n209 ;
  assign n211 = ioin114 & n205 ;
  assign n212 = n210 | n211 ;
  assign n213 = n206 & n212 ;
  assign n214 = ioin115 | n213 ;
  assign n215 = iofn3 & n89 ;
  assign n216 = ioin215 & n215 ;
  assign n217 = ioin215 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ioin115 & n213 ;
  assign n220 = n218 | n219 ;
  assign n221 = n214 & n220 ;
  assign n222 = ioin116 & n221 ;
  assign n223 = iofn3 & n90 ;
  assign n224 = ~ioin216 & n223 ;
  assign n225 = ioin216 & ~n223 ;
  assign n226 = n224 | n225 ;
  assign n227 = ioin116 | n221 ;
  assign n228 = n226 & n227 ;
  assign n229 = n222 | n228 ;
  assign n230 = ioin117 & n229 ;
  assign n231 = iofn3 & n91 ;
  assign n232 = ioin217 & n231 ;
  assign n233 = ioin217 | n231 ;
  assign n234 = ~n232 & n233 ;
  assign n235 = ioin117 | n229 ;
  assign n236 = n234 & n235 ;
  assign n237 = n230 | n236 ;
  assign n238 = ioin118 & n237 ;
  assign n239 = iofn3 & n92 ;
  assign n240 = ~ioin218 & n239 ;
  assign n241 = ioin218 & ~n239 ;
  assign n242 = n240 | n241 ;
  assign n243 = ioin118 | n237 ;
  assign n244 = n242 & n243 ;
  assign n245 = n238 | n244 ;
  assign n246 = ioin119 | n245 ;
  assign n247 = iofn3 & n93 ;
  assign n248 = ioin219 & n247 ;
  assign n249 = ioin219 | n247 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = ioin119 & n245 ;
  assign n252 = n250 | n251 ;
  assign n253 = n246 & n252 ;
  assign n254 = ioin120 | n253 ;
  assign n255 = iofn3 & n94 ;
  assign n256 = ~ioin220 & n255 ;
  assign n257 = ioin220 & ~n255 ;
  assign n258 = n256 | n257 ;
  assign n259 = ioin120 & n253 ;
  assign n260 = n258 | n259 ;
  assign n261 = n254 & n260 ;
  assign n262 = ioin121 | n261 ;
  assign n263 = iofn3 & n95 ;
  assign n264 = ioin221 & n263 ;
  assign n265 = ioin221 | n263 ;
  assign n266 = ~n264 & n265 ;
  assign n267 = ioin121 & n261 ;
  assign n268 = n266 | n267 ;
  assign n269 = n262 & n268 ;
  assign n270 = ioin122 & n269 ;
  assign n271 = ioin122 | n269 ;
  assign n272 = ~n270 & n271 ;
  assign n273 = n100 | n272 ;
  assign n274 = n100 & n272 ;
  assign n275 = n273 & ~n274 ;
  assign n276 = ~n75 & n275 ;
  assign n277 = iofn0 & ~iofn1 ;
  assign n278 = iofn2 & ~iofn3 ;
  assign n279 = n277 & n278 ;
  assign n280 = ~iofn2 & iofn3 ;
  assign n281 = iofn0 & iofn1 ;
  assign n282 = n280 & n281 ;
  assign n283 = n279 | n282 ;
  assign n284 = ~iofn0 & n278 ;
  assign n285 = ioin122 | n284 ;
  assign n286 = ioin222 & n285 ;
  assign n287 = n278 & n281 ;
  assign n288 = ioin122 & ~n287 ;
  assign n289 = n286 | n288 ;
  assign n290 = ~n72 & n277 ;
  assign n291 = ~n73 & n278 ;
  assign n292 = ioin222 & n291 ;
  assign n293 = n288 & n292 ;
  assign n294 = n290 | n293 ;
  assign n295 = n289 & ~n294 ;
  assign n296 = n283 | n295 ;
  assign n297 = ioin116 & ~n283 ;
  assign n298 = ioin115 & n283 ;
  assign n299 = n297 | n298 ;
  assign n300 = ioin20 | n299 ;
  assign n301 = ioin115 & ~n283 ;
  assign n302 = ioin116 & n283 ;
  assign n303 = n301 | n302 ;
  assign n304 = ioin20 & ~n303 ;
  assign n305 = n300 & ~n304 ;
  assign n306 = ioin21 & n305 ;
  assign n307 = ioin114 & n283 ;
  assign n308 = ioin117 & ~n283 ;
  assign n309 = n307 | n308 ;
  assign n310 = ioin20 & n309 ;
  assign n311 = ioin118 & ~n283 ;
  assign n312 = ioin113 & n283 ;
  assign n313 = n311 | n312 ;
  assign n314 = ~ioin20 & n313 ;
  assign n315 = n310 | n314 ;
  assign n316 = ~ioin21 & n315 ;
  assign n317 = n306 | n316 ;
  assign n318 = ioin22 & n317 ;
  assign n319 = ioin112 & n283 ;
  assign n320 = ioin119 & ~n283 ;
  assign n321 = n319 | n320 ;
  assign n322 = ioin20 & n321 ;
  assign n323 = ioin111 & n283 ;
  assign n324 = ioin120 & ~n283 ;
  assign n325 = n323 | n324 ;
  assign n326 = ~ioin20 & n325 ;
  assign n327 = n322 | n326 ;
  assign n328 = ioin21 & n327 ;
  assign n329 = ioin110 & n283 ;
  assign n330 = ioin121 & ~n283 ;
  assign n331 = n329 | n330 ;
  assign n332 = ioin20 & n331 ;
  assign n333 = ioin19 & n283 ;
  assign n334 = ioin122 & ~n283 ;
  assign n335 = n333 | n334 ;
  assign n336 = ~ioin20 & n335 ;
  assign n337 = n332 | n336 ;
  assign n338 = ~ioin21 & n337 ;
  assign n339 = n328 | n338 ;
  assign n340 = ~ioin22 & n339 ;
  assign n341 = n318 | n340 ;
  assign n342 = ~ioin23 & n341 ;
  assign n343 = ioin114 & ~n283 ;
  assign n344 = ioin117 & n283 ;
  assign n345 = n343 | n344 ;
  assign n346 = ~ioin20 & n345 ;
  assign n347 = ioin113 & ~n283 ;
  assign n348 = ioin118 & n283 ;
  assign n349 = n347 | n348 ;
  assign n350 = ioin20 & n349 ;
  assign n351 = n346 | n350 ;
  assign n352 = ~ioin21 & n351 ;
  assign n353 = ioin112 & ~n283 ;
  assign n354 = ioin119 & n283 ;
  assign n355 = n353 | n354 ;
  assign n356 = ~ioin20 & n355 ;
  assign n357 = ioin111 & ~n283 ;
  assign n358 = ioin120 & n283 ;
  assign n359 = n357 | n358 ;
  assign n360 = ioin20 & n359 ;
  assign n361 = n356 | n360 ;
  assign n362 = ioin21 & n361 ;
  assign n363 = n352 | n362 ;
  assign n364 = ~ioin22 & n363 ;
  assign n365 = ioin110 & ~n283 ;
  assign n366 = ioin121 & n283 ;
  assign n367 = n365 | n366 ;
  assign n368 = ~ioin20 & n367 ;
  assign n369 = ioin19 & ~n283 ;
  assign n370 = ioin122 & n283 ;
  assign n371 = n369 | n370 ;
  assign n372 = ioin20 & n371 ;
  assign n373 = n368 | n372 ;
  assign n374 = ~ioin21 & n373 ;
  assign n375 = ioin17 & ~n283 ;
  assign n376 = ioin124 & n283 ;
  assign n377 = n375 | n376 ;
  assign n378 = ioin20 & n377 ;
  assign n379 = ioin123 & n283 ;
  assign n380 = ioin18 & ~n283 ;
  assign n381 = n379 | n380 ;
  assign n382 = ~ioin20 & n381 ;
  assign n383 = n378 | n382 ;
  assign n384 = ioin21 & n383 ;
  assign n385 = n374 | n384 ;
  assign n386 = ioin22 & n385 ;
  assign n387 = n364 | n386 ;
  assign n388 = ioin23 & n387 ;
  assign n389 = ioin24 | n388 ;
  assign n390 = n342 | n389 ;
  assign n391 = ioin10 & ~n283 ;
  assign n392 = ioin131 & n283 ;
  assign n393 = n391 | n392 ;
  assign n394 = iofn3 & n393 ;
  assign n395 = ioin23 & n394 ;
  assign n396 = ioin125 & n283 ;
  assign n397 = ioin16 & ~n283 ;
  assign n398 = n396 | n397 ;
  assign n399 = ~ioin20 & n398 ;
  assign n400 = ioin15 & ~n283 ;
  assign n401 = ioin126 & n283 ;
  assign n402 = n400 | n401 ;
  assign n403 = ioin20 & n402 ;
  assign n404 = n399 | n403 ;
  assign n405 = ~ioin21 & n404 ;
  assign n406 = ioin14 & ~n283 ;
  assign n407 = ioin127 & n283 ;
  assign n408 = n406 | n407 ;
  assign n409 = ~ioin20 & n408 ;
  assign n410 = ioin13 & ~n283 ;
  assign n411 = ioin128 & n283 ;
  assign n412 = n410 | n411 ;
  assign n413 = ioin20 & n412 ;
  assign n414 = n409 | n413 ;
  assign n415 = ioin21 & n414 ;
  assign n416 = n405 | n415 ;
  assign n417 = ~ioin22 & n416 ;
  assign n418 = ioin12 & ~n283 ;
  assign n419 = ioin129 & n283 ;
  assign n420 = n418 | n419 ;
  assign n421 = ~ioin20 & n420 ;
  assign n422 = ioin11 & ~n283 ;
  assign n423 = ioin130 & n283 ;
  assign n424 = n422 | n423 ;
  assign n425 = ioin20 & n424 ;
  assign n426 = n421 | n425 ;
  assign n427 = ioin21 | n426 ;
  assign n428 = ioin21 & ~n394 ;
  assign n429 = ~ioin20 & n393 ;
  assign n430 = n428 & ~n429 ;
  assign n431 = n427 & ~n430 ;
  assign n432 = ioin22 & n431 ;
  assign n433 = n417 | n432 ;
  assign n434 = ~ioin23 & n433 ;
  assign n435 = n395 | n434 ;
  assign n436 = ioin24 & ~n435 ;
  assign n437 = n390 & ~n436 ;
  assign n438 = n290 & n437 ;
  assign n439 = n296 | n438 ;
  assign n440 = iofn2 & n69 ;
  assign n441 = n75 & ~n440 ;
  assign n442 = ioin24 & n394 ;
  assign n443 = ~ioin20 & n371 ;
  assign n444 = ioin20 & n381 ;
  assign n445 = n443 | n444 ;
  assign n446 = ~ioin21 & n445 ;
  assign n447 = ~ioin20 & n377 ;
  assign n448 = ioin20 & n398 ;
  assign n449 = n447 | n448 ;
  assign n450 = ioin21 & n449 ;
  assign n451 = n446 | n450 ;
  assign n452 = ~ioin22 & n451 ;
  assign n453 = ~ioin20 & n402 ;
  assign n454 = ioin20 & n408 ;
  assign n455 = n453 | n454 ;
  assign n456 = ~ioin21 & n455 ;
  assign n457 = ~ioin20 & n412 ;
  assign n458 = ioin20 & n420 ;
  assign n459 = n457 | n458 ;
  assign n460 = ioin21 & n459 ;
  assign n461 = n456 | n460 ;
  assign n462 = ioin22 & n461 ;
  assign n463 = n452 | n462 ;
  assign n464 = ioin23 | n463 ;
  assign n465 = ioin22 & n394 ;
  assign n466 = ~ioin20 & n424 ;
  assign n467 = ioin20 & n393 ;
  assign n468 = n466 | n467 ;
  assign n469 = ioin21 | n468 ;
  assign n470 = ~n428 & n469 ;
  assign n471 = ~ioin22 & n470 ;
  assign n472 = n465 | n471 ;
  assign n473 = ioin23 & ~n472 ;
  assign n474 = n464 & ~n473 ;
  assign n475 = ~ioin24 & n474 ;
  assign n476 = n442 | n475 ;
  assign n477 = n283 & ~n476 ;
  assign n478 = n441 & ~n477 ;
  assign n479 = n439 & n478 ;
  assign n480 = n276 | n479 ;
  assign n481 = n150 & ~n151 ;
  assign n482 = ~n155 & n481 ;
  assign n483 = n155 & ~n481 ;
  assign n484 = n482 | n483 ;
  assign n485 = ~n75 & n484 ;
  assign n486 = ~ioin21 & n305 ;
  assign n487 = ioin21 & n351 ;
  assign n488 = n486 | n487 ;
  assign n489 = ~ioin22 & n488 ;
  assign n490 = ~ioin21 & n361 ;
  assign n491 = ioin21 & n373 ;
  assign n492 = n490 | n491 ;
  assign n493 = ioin22 & n492 ;
  assign n494 = n489 | n493 ;
  assign n495 = ioin23 & n494 ;
  assign n496 = ioin21 & n315 ;
  assign n497 = ~ioin21 & n327 ;
  assign n498 = n496 | n497 ;
  assign n499 = ioin22 & n498 ;
  assign n500 = ioin21 & n337 ;
  assign n501 = ioin17 & n283 ;
  assign n502 = ioin124 & ~n283 ;
  assign n503 = n501 | n502 ;
  assign n504 = ~ioin20 & n503 ;
  assign n505 = ioin123 & ~n283 ;
  assign n506 = ioin18 & n283 ;
  assign n507 = n505 | n506 ;
  assign n508 = ioin20 & n507 ;
  assign n509 = n504 | n508 ;
  assign n510 = ~ioin21 & n509 ;
  assign n511 = n500 | n510 ;
  assign n512 = ~ioin22 & n511 ;
  assign n513 = n499 | n512 ;
  assign n514 = ~ioin23 & n513 ;
  assign n515 = n495 | n514 ;
  assign n516 = ioin24 | n515 ;
  assign n517 = ~ioin21 & n383 ;
  assign n518 = ioin21 & n404 ;
  assign n519 = n517 | n518 ;
  assign n520 = ~ioin22 & n519 ;
  assign n521 = ~ioin21 & n414 ;
  assign n522 = ioin21 & n426 ;
  assign n523 = n521 | n522 ;
  assign n524 = ioin22 & n523 ;
  assign n525 = n520 | n524 ;
  assign n526 = ~ioin23 & n525 ;
  assign n527 = ~iofn3 & n77 ;
  assign n528 = ioin23 & ~n527 ;
  assign n529 = n393 & n528 ;
  assign n530 = n526 | n529 ;
  assign n531 = ioin24 & ~n530 ;
  assign n532 = n516 & ~n531 ;
  assign n533 = n283 & ~n532 ;
  assign n534 = n441 & ~n533 ;
  assign n535 = ioin17 & ~n287 ;
  assign n536 = ioin27 & n291 ;
  assign n537 = n535 & n536 ;
  assign n538 = n290 | n537 ;
  assign n539 = ioin17 | n284 ;
  assign n540 = ioin27 & n539 ;
  assign n541 = n535 | n540 ;
  assign n542 = ~n538 & n541 ;
  assign n543 = n283 | n542 ;
  assign n544 = ~ioin21 & n449 ;
  assign n545 = ioin21 & n455 ;
  assign n546 = n544 | n545 ;
  assign n547 = ~ioin22 & n546 ;
  assign n548 = ~ioin21 & n459 ;
  assign n549 = ioin21 & n468 ;
  assign n550 = n548 | n549 ;
  assign n551 = ioin22 & n550 ;
  assign n552 = n547 | n551 ;
  assign n553 = ~ioin23 & n552 ;
  assign n554 = n395 | n553 ;
  assign n555 = ~ioin24 & n554 ;
  assign n556 = n442 | n555 ;
  assign n557 = n290 & n556 ;
  assign n558 = n543 | n557 ;
  assign n559 = n534 & n558 ;
  assign n560 = n485 | n559 ;
  assign n561 = ioin222 | n96 ;
  assign n562 = ioin223 | n561 ;
  assign n563 = ioin224 | n562 ;
  assign n564 = ioin225 | n563 ;
  assign n565 = ioin226 | n564 ;
  assign n566 = ioin227 | n565 ;
  assign n567 = iofn3 & n566 ;
  assign n568 = ioin228 | n567 ;
  assign n569 = iofn3 & n568 ;
  assign n570 = ioin229 | n569 ;
  assign n571 = iofn3 & n570 ;
  assign n572 = ioin230 & iofn3 ;
  assign n573 = n571 | n572 ;
  assign n574 = ~ioin231 & n573 ;
  assign n575 = ioin231 & ~n573 ;
  assign n576 = n574 | n575 ;
  assign n577 = ioin131 | n576 ;
  assign n578 = ioin131 & n576 ;
  assign n579 = iofn3 & n565 ;
  assign n580 = ~ioin227 & n579 ;
  assign n581 = ioin227 & ~n579 ;
  assign n582 = n580 | n581 ;
  assign n583 = n100 & n271 ;
  assign n584 = n270 | n583 ;
  assign n585 = ioin123 | n584 ;
  assign n586 = iofn3 & n561 ;
  assign n587 = ioin223 & n586 ;
  assign n588 = ioin223 | n586 ;
  assign n589 = ~n587 & n588 ;
  assign n590 = ioin123 & n584 ;
  assign n591 = n589 | n590 ;
  assign n592 = n585 & n591 ;
  assign n593 = ioin124 & n592 ;
  assign n594 = iofn3 & n562 ;
  assign n595 = ~ioin224 & n594 ;
  assign n596 = ioin224 & ~n594 ;
  assign n597 = n595 | n596 ;
  assign n598 = ioin124 | n592 ;
  assign n599 = n597 & n598 ;
  assign n600 = n593 | n599 ;
  assign n601 = ioin125 & n600 ;
  assign n602 = iofn3 & n563 ;
  assign n603 = ioin225 & ~n602 ;
  assign n604 = ~ioin225 & n602 ;
  assign n605 = n603 | n604 ;
  assign n606 = ioin125 | n600 ;
  assign n607 = n605 & n606 ;
  assign n608 = n601 | n607 ;
  assign n609 = ioin126 & n608 ;
  assign n610 = iofn3 & n564 ;
  assign n611 = ioin226 & n610 ;
  assign n612 = ioin226 | n610 ;
  assign n613 = ~n611 & n612 ;
  assign n614 = ioin126 | n608 ;
  assign n615 = n613 & n614 ;
  assign n616 = n609 | n615 ;
  assign n617 = ioin127 & n616 ;
  assign n618 = n582 | n617 ;
  assign n619 = ioin127 | n616 ;
  assign n620 = n618 & n619 ;
  assign n621 = ioin128 & n620 ;
  assign n622 = ioin228 & n567 ;
  assign n623 = n568 & ~n622 ;
  assign n624 = ioin128 | n620 ;
  assign n625 = n623 & n624 ;
  assign n626 = n621 | n625 ;
  assign n627 = ioin129 | n626 ;
  assign n628 = ioin229 & n569 ;
  assign n629 = n570 & ~n628 ;
  assign n630 = ioin129 & n626 ;
  assign n631 = n629 | n630 ;
  assign n632 = n627 & n631 ;
  assign n633 = ioin130 & n632 ;
  assign n634 = ioin230 & n571 ;
  assign n635 = ioin230 | n571 ;
  assign n636 = ~n634 & n635 ;
  assign n637 = ioin130 | n632 ;
  assign n638 = n636 & n637 ;
  assign n639 = n633 | n638 ;
  assign n640 = n578 | n639 ;
  assign n641 = n577 & n640 ;
  assign n642 = ~n230 & n235 ;
  assign n643 = ~n234 & n642 ;
  assign n644 = n234 & ~n642 ;
  assign n645 = n643 | n644 ;
  assign n646 = ~n609 & n614 ;
  assign n647 = ~n613 & n646 ;
  assign n648 = n613 & ~n646 ;
  assign n649 = n647 | n648 ;
  assign n650 = n102 & ~n103 ;
  assign n651 = n108 | n650 ;
  assign n652 = n108 & n650 ;
  assign n653 = n651 & ~n652 ;
  assign n654 = n585 & ~n590 ;
  assign n655 = ~n589 & n654 ;
  assign n656 = n589 & ~n654 ;
  assign n657 = n655 | n656 ;
  assign n658 = ~n75 & n653 ;
  assign n659 = ioin23 & n341 ;
  assign n660 = ioin130 & ~n283 ;
  assign n661 = ioin11 & n283 ;
  assign n662 = n660 | n661 ;
  assign n663 = ~n76 & n662 ;
  assign n664 = ioin22 | n663 ;
  assign n665 = ~ioin21 & ioin20 ;
  assign n666 = ioin129 & ~n283 ;
  assign n667 = ioin12 & n283 ;
  assign n668 = n666 | n667 ;
  assign n669 = n665 & n668 ;
  assign n670 = n664 | n669 ;
  assign n671 = ioin128 & ~n283 ;
  assign n672 = ioin13 & n283 ;
  assign n673 = n671 | n672 ;
  assign n674 = ~ioin20 & n673 ;
  assign n675 = ioin127 & ~n283 ;
  assign n676 = ioin14 & n283 ;
  assign n677 = n675 | n676 ;
  assign n678 = ioin20 & n677 ;
  assign n679 = n674 | n678 ;
  assign n680 = ioin21 & n679 ;
  assign n681 = n670 | n680 ;
  assign n682 = ioin126 & ~n283 ;
  assign n683 = ioin15 & n283 ;
  assign n684 = n682 | n683 ;
  assign n685 = ~ioin20 & n684 ;
  assign n686 = ioin125 & ~n283 ;
  assign n687 = ioin16 & n283 ;
  assign n688 = n686 | n687 ;
  assign n689 = ioin20 & n688 ;
  assign n690 = n685 | n689 ;
  assign n691 = ~ioin21 & n690 ;
  assign n692 = ioin21 & n509 ;
  assign n693 = n691 | n692 ;
  assign n694 = ioin22 & ~n693 ;
  assign n695 = n681 & ~n694 ;
  assign n696 = ~ioin23 & n695 ;
  assign n697 = n659 | n696 ;
  assign n698 = ~ioin24 & n697 ;
  assign n699 = ~ioin23 & n387 ;
  assign n700 = ioin23 & n433 ;
  assign n701 = n699 | n700 ;
  assign n702 = ioin24 & n701 ;
  assign n703 = n698 | n702 ;
  assign n704 = n283 & ~n703 ;
  assign n705 = n441 & ~n704 ;
  assign n706 = ioin21 & ioin11 ;
  assign n707 = n287 & ~n706 ;
  assign n708 = n290 | n707 ;
  assign n709 = ioin21 & n284 ;
  assign n710 = ioin11 | n709 ;
  assign n711 = n291 & n706 ;
  assign n712 = n710 & ~n711 ;
  assign n713 = n287 | n712 ;
  assign n714 = ~n708 & n713 ;
  assign n715 = n283 | n714 ;
  assign n716 = ~ioin23 & n472 ;
  assign n717 = n395 | n716 ;
  assign n718 = ~ioin24 & n717 ;
  assign n719 = n442 | n718 ;
  assign n720 = n290 & n719 ;
  assign n721 = n715 | n720 ;
  assign n722 = n705 & n721 ;
  assign n723 = n658 | n722 ;
  assign n724 = n158 & ~n159 ;
  assign n725 = n163 | n724 ;
  assign n726 = n163 & n724 ;
  assign n727 = n725 & ~n726 ;
  assign n728 = ioin10 | ioin20 ;
  assign n729 = ~n101 & n728 ;
  assign n730 = n214 & ~n219 ;
  assign n731 = n218 & ~n730 ;
  assign n732 = ~n218 & n730 ;
  assign n733 = n731 | n732 ;
  assign n734 = ~n75 & n733 ;
  assign n735 = ioin23 | n494 ;
  assign n736 = ~ioin24 & n735 ;
  assign n737 = ioin23 & ~n525 ;
  assign n738 = n736 & ~n737 ;
  assign n739 = ~iofn3 & n78 ;
  assign n740 = ioin24 & ~n739 ;
  assign n741 = n393 & n740 ;
  assign n742 = n738 | n741 ;
  assign n743 = n283 & ~n742 ;
  assign n744 = n441 & ~n743 ;
  assign n745 = ioin115 | n284 ;
  assign n746 = ioin115 & ~n287 ;
  assign n747 = ioin215 & ~n746 ;
  assign n748 = n745 & n747 ;
  assign n749 = ioin215 & n291 ;
  assign n750 = n746 & ~n749 ;
  assign n751 = n748 | n750 ;
  assign n752 = ~n290 & n751 ;
  assign n753 = n283 | n752 ;
  assign n754 = ~ioin20 & n303 ;
  assign n755 = ioin20 & n345 ;
  assign n756 = n754 | n755 ;
  assign n757 = ~ioin21 & n756 ;
  assign n758 = ~ioin20 & n349 ;
  assign n759 = ioin20 & n355 ;
  assign n760 = n758 | n759 ;
  assign n761 = ioin21 & n760 ;
  assign n762 = n757 | n761 ;
  assign n763 = ~ioin22 & n762 ;
  assign n764 = ~ioin20 & n359 ;
  assign n765 = ioin20 & n367 ;
  assign n766 = n764 | n765 ;
  assign n767 = ~ioin21 & n766 ;
  assign n768 = ioin21 & n445 ;
  assign n769 = n767 | n768 ;
  assign n770 = ioin22 & n769 ;
  assign n771 = n763 | n770 ;
  assign n772 = ~ioin23 & n771 ;
  assign n773 = ioin23 & n552 ;
  assign n774 = n772 | n773 ;
  assign n775 = ~ioin24 & n774 ;
  assign n776 = n442 | n775 ;
  assign n777 = n290 & n776 ;
  assign n778 = n753 | n777 ;
  assign n779 = n744 & n778 ;
  assign n780 = n734 | n779 ;
  assign n781 = n577 & ~n578 ;
  assign n782 = n639 & ~n781 ;
  assign n783 = ~n639 & n781 ;
  assign n784 = n782 | n783 ;
  assign n785 = ~n75 & n784 ;
  assign n786 = ~iofn3 & n79 ;
  assign n787 = n393 & ~n786 ;
  assign n788 = n283 & ~n787 ;
  assign n789 = n441 & ~n788 ;
  assign n790 = ioin131 & ioin231 ;
  assign n791 = n287 & ~n790 ;
  assign n792 = n290 | n791 ;
  assign n793 = ioin131 & ~n291 ;
  assign n794 = ~ioin131 & ioin231 ;
  assign n795 = n284 & n794 ;
  assign n796 = ioin131 & ~ioin231 ;
  assign n797 = n795 | n796 ;
  assign n798 = n793 | n797 ;
  assign n799 = ~n792 & n798 ;
  assign n800 = n283 | n799 ;
  assign n801 = n662 & n665 ;
  assign n802 = ~ioin20 & n668 ;
  assign n803 = ioin20 & n673 ;
  assign n804 = n802 | n803 ;
  assign n805 = ioin21 & n804 ;
  assign n806 = n801 | n805 ;
  assign n807 = ioin131 | n283 ;
  assign n808 = ~n76 & n807 ;
  assign n809 = ~ioin10 & n283 ;
  assign n810 = n808 & ~n809 ;
  assign n811 = ioin22 | n810 ;
  assign n812 = n806 | n811 ;
  assign n813 = ~ioin20 & n677 ;
  assign n814 = ioin20 & n684 ;
  assign n815 = n813 | n814 ;
  assign n816 = ~ioin21 & n815 ;
  assign n817 = ioin20 & n503 ;
  assign n818 = ~ioin20 & n688 ;
  assign n819 = n817 | n818 ;
  assign n820 = ioin21 & n819 ;
  assign n821 = n816 | n820 ;
  assign n822 = ioin22 & ~n821 ;
  assign n823 = n812 & ~n822 ;
  assign n824 = ~ioin23 & n823 ;
  assign n825 = ioin20 & n299 ;
  assign n826 = ~ioin20 & n309 ;
  assign n827 = n825 | n826 ;
  assign n828 = ioin21 & n827 ;
  assign n829 = ioin20 & n313 ;
  assign n830 = ~ioin20 & n321 ;
  assign n831 = n829 | n830 ;
  assign n832 = ~ioin21 & n831 ;
  assign n833 = n828 | n832 ;
  assign n834 = ioin22 & n833 ;
  assign n835 = ioin20 & n325 ;
  assign n836 = ~ioin20 & n331 ;
  assign n837 = n835 | n836 ;
  assign n838 = ioin21 & n837 ;
  assign n839 = ioin20 & n335 ;
  assign n840 = ~ioin20 & n507 ;
  assign n841 = n839 | n840 ;
  assign n842 = ~ioin21 & n841 ;
  assign n843 = n838 | n842 ;
  assign n844 = ~ioin22 & n843 ;
  assign n845 = n834 | n844 ;
  assign n846 = ioin23 & n845 ;
  assign n847 = n824 | n846 ;
  assign n848 = ~ioin24 & n847 ;
  assign n849 = ioin24 & n774 ;
  assign n850 = n848 | n849 ;
  assign n851 = n290 & n850 ;
  assign n852 = n800 | n851 ;
  assign n853 = n789 & n852 ;
  assign n854 = n785 | n853 ;
  assign n855 = n174 & ~n179 ;
  assign n856 = n178 | n855 ;
  assign n857 = n178 & n855 ;
  assign n858 = n856 & ~n857 ;
  assign n859 = ~n601 & n606 ;
  assign n860 = n605 | n859 ;
  assign n861 = n605 & n859 ;
  assign n862 = n860 & ~n861 ;
  assign n863 = ~n75 & n862 ;
  assign n864 = ~ioin24 & n435 ;
  assign n865 = n442 | n864 ;
  assign n866 = n283 & ~n865 ;
  assign n867 = n441 & ~n866 ;
  assign n868 = ioin225 & ioin125 ;
  assign n869 = n287 & ~n868 ;
  assign n870 = n290 | n869 ;
  assign n871 = ioin225 & n284 ;
  assign n872 = ioin125 | n871 ;
  assign n873 = n291 & n868 ;
  assign n874 = n872 & ~n873 ;
  assign n875 = n287 | n874 ;
  assign n876 = ~n870 & n875 ;
  assign n877 = n283 | n876 ;
  assign n878 = ~ioin21 & n827 ;
  assign n879 = ioin21 & n756 ;
  assign n880 = n878 | n879 ;
  assign n881 = ~ioin22 & n880 ;
  assign n882 = ~ioin21 & n760 ;
  assign n883 = ioin21 & n766 ;
  assign n884 = n882 | n883 ;
  assign n885 = ioin22 & n884 ;
  assign n886 = n881 | n885 ;
  assign n887 = ioin23 & ~n886 ;
  assign n888 = ioin21 & n831 ;
  assign n889 = ~ioin21 & n837 ;
  assign n890 = n888 | n889 ;
  assign n891 = ioin22 & ~n890 ;
  assign n892 = ~ioin21 & n819 ;
  assign n893 = ioin21 & n841 ;
  assign n894 = n892 | n893 ;
  assign n895 = ioin22 | n894 ;
  assign n896 = ~n891 & n895 ;
  assign n897 = ioin23 | n896 ;
  assign n898 = ~n887 & n897 ;
  assign n899 = ~ioin24 & n898 ;
  assign n900 = ioin24 & n474 ;
  assign n901 = n899 | n900 ;
  assign n902 = n290 & n901 ;
  assign n903 = n877 | n902 ;
  assign n904 = n867 & n903 ;
  assign n905 = n863 | n904 ;
  assign n906 = ~n75 & n858 ;
  assign n907 = ioin110 | n284 ;
  assign n908 = ioin110 & ~n287 ;
  assign n909 = ioin210 & ~n908 ;
  assign n910 = n907 & n909 ;
  assign n911 = ioin210 & n291 ;
  assign n912 = n908 & ~n911 ;
  assign n913 = n910 | n912 ;
  assign n914 = ~n290 & n913 ;
  assign n915 = n283 | n914 ;
  assign n916 = ~ioin22 & n385 ;
  assign n917 = ioin22 & n416 ;
  assign n918 = n916 | n917 ;
  assign n919 = ioin23 | n918 ;
  assign n920 = ~ioin22 & n431 ;
  assign n921 = n465 | n920 ;
  assign n922 = ioin23 & ~n921 ;
  assign n923 = n919 & ~n922 ;
  assign n924 = ~ioin24 & n923 ;
  assign n925 = n442 | n924 ;
  assign n926 = n290 & n925 ;
  assign n927 = n915 | n926 ;
  assign n928 = ioin22 & n880 ;
  assign n929 = ~ioin22 & n890 ;
  assign n930 = n928 | n929 ;
  assign n931 = ~ioin23 & n930 ;
  assign n932 = ~ioin22 & n884 ;
  assign n933 = ioin22 & n451 ;
  assign n934 = n932 | n933 ;
  assign n935 = ioin23 & n934 ;
  assign n936 = ioin24 | n935 ;
  assign n937 = n931 | n936 ;
  assign n938 = ioin22 | n461 ;
  assign n939 = ioin22 & ~n470 ;
  assign n940 = n938 & ~n939 ;
  assign n941 = ~ioin23 & n940 ;
  assign n942 = n395 | n941 ;
  assign n943 = ioin24 & ~n942 ;
  assign n944 = n937 & ~n943 ;
  assign n945 = n283 & ~n944 ;
  assign n946 = n441 & ~n945 ;
  assign n947 = n927 & n946 ;
  assign n948 = n906 | n947 ;
  assign n949 = n206 & ~n211 ;
  assign n950 = n210 & n949 ;
  assign n951 = n210 | n949 ;
  assign n952 = ~n950 & n951 ;
  assign n953 = ~n75 & n952 ;
  assign n954 = ioin214 & ioin114 ;
  assign n955 = n287 & ~n954 ;
  assign n956 = n290 | n955 ;
  assign n957 = ioin214 & n284 ;
  assign n958 = ioin114 | n957 ;
  assign n959 = n291 & n954 ;
  assign n960 = n958 & ~n959 ;
  assign n961 = n287 | n960 ;
  assign n962 = ~n956 & n961 ;
  assign n963 = n283 | n962 ;
  assign n964 = ~ioin24 & n701 ;
  assign n965 = n442 | n964 ;
  assign n966 = n290 & n965 ;
  assign n967 = n963 | n966 ;
  assign n968 = ioin23 | n886 ;
  assign n969 = ioin23 & ~n463 ;
  assign n970 = n968 & ~n969 ;
  assign n971 = ~ioin24 & n970 ;
  assign n972 = ioin24 & n717 ;
  assign n973 = n971 | n972 ;
  assign n974 = n283 & ~n973 ;
  assign n975 = n441 & ~n974 ;
  assign n976 = n967 & n975 ;
  assign n977 = n953 | n976 ;
  assign n978 = ~n593 & n598 ;
  assign n979 = n597 | n978 ;
  assign n980 = n597 & n978 ;
  assign n981 = n979 & ~n980 ;
  assign n982 = ~n75 & n981 ;
  assign n983 = ioin224 & ioin124 ;
  assign n984 = n287 & ~n983 ;
  assign n985 = n290 | n984 ;
  assign n986 = ioin224 & n284 ;
  assign n987 = ioin124 | n986 ;
  assign n988 = n291 & n983 ;
  assign n989 = n987 & ~n988 ;
  assign n990 = n287 | n989 ;
  assign n991 = ~n985 & n990 ;
  assign n992 = n283 | n991 ;
  assign n993 = n290 & n532 ;
  assign n994 = n992 | n993 ;
  assign n995 = n283 & ~n556 ;
  assign n996 = n441 & ~n995 ;
  assign n997 = n994 & n996 ;
  assign n998 = n982 | n997 ;
  assign n999 = n134 & ~n135 ;
  assign n1000 = n139 & ~n999 ;
  assign n1001 = ~n139 & n999 ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = n190 & ~n195 ;
  assign n1004 = n194 & n1003 ;
  assign n1005 = n194 | n1003 ;
  assign n1006 = ~n1004 & n1005 ;
  assign n1007 = ~n75 & n1006 ;
  assign n1008 = ioin112 | n284 ;
  assign n1009 = ioin212 & n1008 ;
  assign n1010 = ioin112 & ~n287 ;
  assign n1011 = n1009 | n1010 ;
  assign n1012 = ioin212 & n291 ;
  assign n1013 = n1010 & n1012 ;
  assign n1014 = n290 | n1013 ;
  assign n1015 = n1011 & ~n1014 ;
  assign n1016 = n283 | n1015 ;
  assign n1017 = ~ioin22 & n492 ;
  assign n1018 = ioin22 & n519 ;
  assign n1019 = n1017 | n1018 ;
  assign n1020 = ~ioin23 & n1019 ;
  assign n1021 = ioin22 | n523 ;
  assign n1022 = ~iofn3 & n76 ;
  assign n1023 = n393 & ~n1022 ;
  assign n1024 = ioin22 & ~n1023 ;
  assign n1025 = n1021 & ~n1024 ;
  assign n1026 = ioin23 & n1025 ;
  assign n1027 = n1020 | n1026 ;
  assign n1028 = ~ioin24 & n1027 ;
  assign n1029 = n442 | n1028 ;
  assign n1030 = n290 & n1029 ;
  assign n1031 = n1016 | n1030 ;
  assign n1032 = ~ioin22 & n833 ;
  assign n1033 = ioin22 & n762 ;
  assign n1034 = n1032 | n1033 ;
  assign n1035 = ioin23 | n1034 ;
  assign n1036 = ~ioin22 & n769 ;
  assign n1037 = ioin22 & n546 ;
  assign n1038 = n1036 | n1037 ;
  assign n1039 = ioin23 & ~n1038 ;
  assign n1040 = n1035 & ~n1039 ;
  assign n1041 = ~ioin24 & n1040 ;
  assign n1042 = ~ioin22 & n550 ;
  assign n1043 = n465 | n1042 ;
  assign n1044 = ~ioin23 & n1043 ;
  assign n1045 = n395 | n1044 ;
  assign n1046 = ioin24 & n1045 ;
  assign n1047 = n1041 | n1046 ;
  assign n1048 = n283 & ~n1047 ;
  assign n1049 = n441 & ~n1048 ;
  assign n1050 = n1031 & n1049 ;
  assign n1051 = n1007 | n1050 ;
  assign n1052 = n166 & ~n171 ;
  assign n1053 = n170 & ~n1052 ;
  assign n1054 = ~n170 & n1052 ;
  assign n1055 = n1053 | n1054 ;
  assign n1056 = ~n633 & n638 ;
  assign n1057 = ~n633 & n637 ;
  assign n1058 = n636 | n1057 ;
  assign n1059 = ~n1056 & n1058 ;
  assign n1060 = n198 & ~n204 ;
  assign n1061 = n198 & ~n203 ;
  assign n1062 = n202 & ~n1061 ;
  assign n1063 = n1060 | n1062 ;
  assign n1064 = ~n75 & n1063 ;
  assign n1065 = ~ioin22 & n317 ;
  assign n1066 = ioin22 & n363 ;
  assign n1067 = n1065 | n1066 ;
  assign n1068 = ioin23 | n1067 ;
  assign n1069 = ioin23 & ~n918 ;
  assign n1070 = n1068 & ~n1069 ;
  assign n1071 = ~ioin24 & n1070 ;
  assign n1072 = ~ioin23 & n921 ;
  assign n1073 = n395 | n1072 ;
  assign n1074 = ioin24 & n1073 ;
  assign n1075 = n1071 | n1074 ;
  assign n1076 = n283 & ~n1075 ;
  assign n1077 = n441 & ~n1076 ;
  assign n1078 = ioin113 | n284 ;
  assign n1079 = ioin213 & n1078 ;
  assign n1080 = ioin113 & ~n287 ;
  assign n1081 = n1079 | n1080 ;
  assign n1082 = ioin213 & n291 ;
  assign n1083 = n1080 & n1082 ;
  assign n1084 = n290 | n1083 ;
  assign n1085 = n1081 & ~n1084 ;
  assign n1086 = n283 | n1085 ;
  assign n1087 = ~ioin23 & n934 ;
  assign n1088 = ioin23 & n940 ;
  assign n1089 = n1087 | n1088 ;
  assign n1090 = ~ioin24 & n1089 ;
  assign n1091 = n442 | n1090 ;
  assign n1092 = n290 & n1091 ;
  assign n1093 = n1086 | n1092 ;
  assign n1094 = n1077 & n1093 ;
  assign n1095 = n1064 | n1094 ;
  assign n1096 = n283 & ~n925 ;
  assign n1097 = n441 & ~n1096 ;
  assign n1098 = ioin221 & ioin121 ;
  assign n1099 = n287 & ~n1098 ;
  assign n1100 = n290 | n1099 ;
  assign n1101 = ioin221 & n284 ;
  assign n1102 = ioin121 | n1101 ;
  assign n1103 = n291 & n1098 ;
  assign n1104 = n1102 & ~n1103 ;
  assign n1105 = n287 | n1104 ;
  assign n1106 = ~n1100 & n1105 ;
  assign n1107 = n283 | n1106 ;
  assign n1108 = n290 & n944 ;
  assign n1109 = n1107 | n1108 ;
  assign n1110 = n1097 & n1109 ;
  assign n1111 = n262 & ~n267 ;
  assign n1112 = n266 & ~n1111 ;
  assign n1113 = ~n266 & n1111 ;
  assign n1114 = n1112 | n1113 ;
  assign n1115 = ~n75 & n1114 ;
  assign n1116 = n1110 | n1115 ;
  assign n1117 = ~n222 & n227 ;
  assign n1118 = n226 | n1117 ;
  assign n1119 = n226 & n1117 ;
  assign n1120 = n1118 & ~n1119 ;
  assign n1121 = ~n75 & n1059 ;
  assign n1122 = ioin130 | n284 ;
  assign n1123 = ioin130 & ~n287 ;
  assign n1124 = ioin230 & ~n1123 ;
  assign n1125 = n1122 & n1124 ;
  assign n1126 = ioin230 & n291 ;
  assign n1127 = n1123 & ~n1126 ;
  assign n1128 = n1125 | n1127 ;
  assign n1129 = ~n290 & n1128 ;
  assign n1130 = n283 | n1129 ;
  assign n1131 = n290 & n703 ;
  assign n1132 = n1130 | n1131 ;
  assign n1133 = n283 & ~n719 ;
  assign n1134 = n441 & ~n1133 ;
  assign n1135 = n1132 & n1134 ;
  assign n1136 = n1121 | n1135 ;
  assign n1137 = n111 & ~n112 ;
  assign n1138 = n115 & ~n1137 ;
  assign n1139 = ~n115 & n1137 ;
  assign n1140 = n1138 | n1139 ;
  assign n1141 = ~n75 & n1140 ;
  assign n1142 = ioin22 & n284 ;
  assign n1143 = ioin12 | n1142 ;
  assign n1144 = ioin12 & ioin22 ;
  assign n1145 = n291 & n1144 ;
  assign n1146 = n1143 & ~n1145 ;
  assign n1147 = n287 | n1146 ;
  assign n1148 = n287 & ~n1144 ;
  assign n1149 = n290 | n1148 ;
  assign n1150 = n1147 & ~n1149 ;
  assign n1151 = n283 | n1150 ;
  assign n1152 = ~ioin24 & n1073 ;
  assign n1153 = n442 | n1152 ;
  assign n1154 = n290 & n1153 ;
  assign n1155 = n1151 | n1154 ;
  assign n1156 = ioin23 & n930 ;
  assign n1157 = ioin24 | n1156 ;
  assign n1158 = ioin22 & ~n894 ;
  assign n1159 = ~ioin21 & n804 ;
  assign n1160 = ioin21 & n815 ;
  assign n1161 = ioin22 | n1160 ;
  assign n1162 = n1159 | n1161 ;
  assign n1163 = ~n1158 & n1162 ;
  assign n1164 = ~ioin23 & n1163 ;
  assign n1165 = n1157 | n1164 ;
  assign n1166 = ioin24 & ~n1089 ;
  assign n1167 = n1165 & ~n1166 ;
  assign n1168 = n283 & ~n1167 ;
  assign n1169 = n441 & ~n1168 ;
  assign n1170 = n1155 & n1169 ;
  assign n1171 = n1141 | n1170 ;
  assign n1172 = ~n75 & n649 ;
  assign n1173 = ioin126 & ~n287 ;
  assign n1174 = ioin126 | n284 ;
  assign n1175 = ioin226 & n1174 ;
  assign n1176 = n1173 | n1175 ;
  assign n1177 = ioin226 & n291 ;
  assign n1178 = n1173 & n1177 ;
  assign n1179 = n290 | n1178 ;
  assign n1180 = n1176 & ~n1179 ;
  assign n1181 = n283 | n1180 ;
  assign n1182 = ioin23 & ~n1067 ;
  assign n1183 = ioin22 & ~n339 ;
  assign n1184 = ioin22 | n693 ;
  assign n1185 = ~n1183 & n1184 ;
  assign n1186 = ioin23 | n1185 ;
  assign n1187 = ~n1182 & n1186 ;
  assign n1188 = ~ioin24 & n1187 ;
  assign n1189 = ioin24 & n923 ;
  assign n1190 = n1188 | n1189 ;
  assign n1191 = n290 & n1190 ;
  assign n1192 = n1181 | n1191 ;
  assign n1193 = ~ioin24 & n942 ;
  assign n1194 = n442 | n1193 ;
  assign n1195 = n283 & ~n1194 ;
  assign n1196 = n441 & ~n1195 ;
  assign n1197 = n1192 & n1196 ;
  assign n1198 = n1172 | n1197 ;
  assign n1199 = ~n75 & n645 ;
  assign n1200 = n283 & ~n965 ;
  assign n1201 = n441 & ~n1200 ;
  assign n1202 = ioin117 & ioin217 ;
  assign n1203 = n287 & ~n1202 ;
  assign n1204 = n290 | n1203 ;
  assign n1205 = ioin217 & n284 ;
  assign n1206 = ioin117 | n1205 ;
  assign n1207 = n291 & n1202 ;
  assign n1208 = n1206 & ~n1207 ;
  assign n1209 = n287 | n1208 ;
  assign n1210 = ~n1204 & n1209 ;
  assign n1211 = n283 | n1210 ;
  assign n1212 = n290 & n973 ;
  assign n1213 = n1211 | n1212 ;
  assign n1214 = n1201 & n1213 ;
  assign n1215 = n1199 | n1214 ;
  assign n1216 = ~n142 & n143 ;
  assign n1217 = n147 | n1216 ;
  assign n1218 = n147 & n1216 ;
  assign n1219 = n1217 & ~n1218 ;
  assign n1220 = ~n238 & n243 ;
  assign n1221 = ~n242 & n1220 ;
  assign n1222 = n242 & ~n1220 ;
  assign n1223 = n1221 | n1222 ;
  assign n1224 = ~n75 & n1223 ;
  assign n1225 = ioin118 & ioin218 ;
  assign n1226 = n287 & ~n1225 ;
  assign n1227 = n290 | n1226 ;
  assign n1228 = ioin218 & n284 ;
  assign n1229 = ioin118 | n1228 ;
  assign n1230 = n291 & n1225 ;
  assign n1231 = n1229 & ~n1230 ;
  assign n1232 = n287 | n1231 ;
  assign n1233 = ~n1227 & n1232 ;
  assign n1234 = n283 | n1233 ;
  assign n1235 = n290 & n1075 ;
  assign n1236 = n1234 | n1235 ;
  assign n1237 = n283 & ~n1091 ;
  assign n1238 = n441 & ~n1237 ;
  assign n1239 = n1236 & n1238 ;
  assign n1240 = n1224 | n1239 ;
  assign n1241 = n75 | n729 ;
  assign n1242 = iofn1 & n440 ;
  assign n1243 = ~n794 & n1242 ;
  assign n1244 = n796 | n1242 ;
  assign n1245 = ~n1243 & n1244 ;
  assign n1246 = n794 | n796 ;
  assign n1247 = n784 & ~n1246 ;
  assign n1248 = n1245 | n1247 ;
  assign n1249 = n440 & n1248 ;
  assign n1250 = n101 & n287 ;
  assign n1251 = ioin10 | n284 ;
  assign n1252 = ~n287 & n728 ;
  assign n1253 = n1251 & n1252 ;
  assign n1254 = n101 & n291 ;
  assign n1255 = n1253 & ~n1254 ;
  assign n1256 = n1250 | n1255 ;
  assign n1257 = ~n290 & n1256 ;
  assign n1258 = n283 | n1257 ;
  assign n1259 = n290 & n787 ;
  assign n1260 = n1258 | n1259 ;
  assign n1261 = ~n440 & n1260 ;
  assign n1262 = n283 & ~n850 ;
  assign n1263 = n1261 & ~n1262 ;
  assign n1264 = n75 & ~n1263 ;
  assign n1265 = ~n1249 & n1264 ;
  assign n1266 = n1241 & ~n1265 ;
  assign n1267 = n126 & ~n127 ;
  assign n1268 = n131 | n1267 ;
  assign n1269 = n131 & n1267 ;
  assign n1270 = n1268 & ~n1269 ;
  assign n1271 = ~n75 & n1270 ;
  assign n1272 = ioin24 & ioin14 ;
  assign n1273 = n287 & ~n1272 ;
  assign n1274 = n290 | n1273 ;
  assign n1275 = ioin24 & n284 ;
  assign n1276 = ioin14 | n1275 ;
  assign n1277 = n291 & n1272 ;
  assign n1278 = n1276 & ~n1277 ;
  assign n1279 = n287 | n1278 ;
  assign n1280 = ~n1274 & n1279 ;
  assign n1281 = n283 | n1280 ;
  assign n1282 = ~ioin23 & n1025 ;
  assign n1283 = n395 | n1282 ;
  assign n1284 = ~ioin24 & n1283 ;
  assign n1285 = n442 | n1284 ;
  assign n1286 = n290 & n1285 ;
  assign n1287 = n1281 | n1286 ;
  assign n1288 = ioin23 & n1034 ;
  assign n1289 = ~ioin22 & n821 ;
  assign n1290 = ioin22 & n843 ;
  assign n1291 = n1289 | n1290 ;
  assign n1292 = ~ioin23 & n1291 ;
  assign n1293 = n1288 | n1292 ;
  assign n1294 = ioin24 | n1293 ;
  assign n1295 = ioin23 | n1038 ;
  assign n1296 = ioin23 & ~n1043 ;
  assign n1297 = n1295 & ~n1296 ;
  assign n1298 = ioin24 & ~n1297 ;
  assign n1299 = n1294 & ~n1298 ;
  assign n1300 = n283 & ~n1299 ;
  assign n1301 = n441 & ~n1300 ;
  assign n1302 = n1287 & n1301 ;
  assign n1303 = n1271 | n1302 ;
  assign n1304 = n246 & ~n251 ;
  assign n1305 = ~n250 & n1304 ;
  assign n1306 = n250 & ~n1304 ;
  assign n1307 = n1305 | n1306 ;
  assign n1308 = ~n75 & n1307 ;
  assign n1309 = n283 & ~n1029 ;
  assign n1310 = n441 & ~n1309 ;
  assign n1311 = ioin219 & n284 ;
  assign n1312 = ioin119 | n1311 ;
  assign n1313 = ioin119 & ioin219 ;
  assign n1314 = n291 & n1313 ;
  assign n1315 = n1312 & ~n1314 ;
  assign n1316 = n287 | n1315 ;
  assign n1317 = n287 & ~n1313 ;
  assign n1318 = n290 | n1317 ;
  assign n1319 = n1316 & ~n1318 ;
  assign n1320 = n283 | n1319 ;
  assign n1321 = n290 & n1047 ;
  assign n1322 = n1320 | n1321 ;
  assign n1323 = n1310 & n1322 ;
  assign n1324 = n1308 | n1323 ;
  assign n1325 = ~n75 & n657 ;
  assign n1326 = ~ioin24 & n530 ;
  assign n1327 = n442 | n1326 ;
  assign n1328 = n283 & ~n1327 ;
  assign n1329 = n441 & ~n1328 ;
  assign n1330 = ioin223 & ioin123 ;
  assign n1331 = n287 & ~n1330 ;
  assign n1332 = n290 | n1331 ;
  assign n1333 = n291 & n1330 ;
  assign n1334 = ioin223 & n284 ;
  assign n1335 = ioin123 | n1334 ;
  assign n1336 = ~n1333 & n1335 ;
  assign n1337 = n287 | n1336 ;
  assign n1338 = ~n1332 & n1337 ;
  assign n1339 = n283 | n1338 ;
  assign n1340 = ioin23 | n845 ;
  assign n1341 = ioin23 & ~n771 ;
  assign n1342 = n1340 & ~n1341 ;
  assign n1343 = ~ioin24 & n1342 ;
  assign n1344 = ioin24 & n554 ;
  assign n1345 = n1343 | n1344 ;
  assign n1346 = n290 & n1345 ;
  assign n1347 = n1339 | n1346 ;
  assign n1348 = n1329 & n1347 ;
  assign n1349 = n1325 | n1348 ;
  assign n1350 = ~n75 & n727 ;
  assign n1351 = ioin18 & ~n287 ;
  assign n1352 = ioin28 & n291 ;
  assign n1353 = n1351 & n1352 ;
  assign n1354 = n290 | n1353 ;
  assign n1355 = ioin18 | n284 ;
  assign n1356 = ioin28 & n1355 ;
  assign n1357 = n1351 | n1356 ;
  assign n1358 = ~n1354 & n1357 ;
  assign n1359 = n283 | n1358 ;
  assign n1360 = n290 & n1327 ;
  assign n1361 = n1359 | n1360 ;
  assign n1362 = n283 & ~n1345 ;
  assign n1363 = n441 & ~n1362 ;
  assign n1364 = n1361 & n1363 ;
  assign n1365 = n1350 | n1364 ;
  assign n1366 = n254 & ~n259 ;
  assign n1367 = n258 | n1366 ;
  assign n1368 = n258 & n1366 ;
  assign n1369 = n1367 & ~n1368 ;
  assign n1370 = ~n75 & n1369 ;
  assign n1371 = ~ioin22 & n498 ;
  assign n1372 = ioin22 & n488 ;
  assign n1373 = n1371 | n1372 ;
  assign n1374 = ~ioin23 & n1373 ;
  assign n1375 = ioin23 & n1019 ;
  assign n1376 = ioin24 | n1375 ;
  assign n1377 = n1374 | n1376 ;
  assign n1378 = ioin24 & ~n1283 ;
  assign n1379 = n1377 & ~n1378 ;
  assign n1380 = n290 & n1379 ;
  assign n1381 = ioin220 & n284 ;
  assign n1382 = ioin120 | n1381 ;
  assign n1383 = ioin120 & ioin220 ;
  assign n1384 = n291 & n1383 ;
  assign n1385 = n1382 & ~n1384 ;
  assign n1386 = n287 | n1385 ;
  assign n1387 = n287 & ~n1383 ;
  assign n1388 = n290 | n1387 ;
  assign n1389 = n1386 & ~n1388 ;
  assign n1390 = n283 | n1389 ;
  assign n1391 = n1380 | n1390 ;
  assign n1392 = ~ioin24 & n1297 ;
  assign n1393 = n442 | n1392 ;
  assign n1394 = n283 & ~n1393 ;
  assign n1395 = n441 & ~n1394 ;
  assign n1396 = n1391 & n1395 ;
  assign n1397 = n1370 | n1396 ;
  assign n1398 = n627 & ~n630 ;
  assign n1399 = n629 & ~n1398 ;
  assign n1400 = ~n629 & n1398 ;
  assign n1401 = n1399 | n1400 ;
  assign n1402 = n118 & ~n119 ;
  assign n1403 = n123 & ~n1402 ;
  assign n1404 = ~n123 & n1402 ;
  assign n1405 = n1403 | n1404 ;
  assign n1406 = ~n75 & n1405 ;
  assign n1407 = ioin23 & n1373 ;
  assign n1408 = ~ioin21 & n679 ;
  assign n1409 = ioin21 & n690 ;
  assign n1410 = n1408 | n1409 ;
  assign n1411 = ~ioin22 & n1410 ;
  assign n1412 = ioin22 & n511 ;
  assign n1413 = n1411 | n1412 ;
  assign n1414 = ~ioin23 & n1413 ;
  assign n1415 = n1407 | n1414 ;
  assign n1416 = ~ioin24 & n1415 ;
  assign n1417 = ioin24 & n1027 ;
  assign n1418 = n1416 | n1417 ;
  assign n1419 = n283 & ~n1418 ;
  assign n1420 = n441 & ~n1419 ;
  assign n1421 = ioin13 & ioin23 ;
  assign n1422 = n287 & n1421 ;
  assign n1423 = ioin23 & n284 ;
  assign n1424 = ioin13 | n1423 ;
  assign n1425 = n291 & n1421 ;
  assign n1426 = n287 | n1425 ;
  assign n1427 = n1424 & ~n1426 ;
  assign n1428 = n1422 | n1427 ;
  assign n1429 = ~n290 & n1428 ;
  assign n1430 = n283 | n1429 ;
  assign n1431 = ~ioin24 & n1045 ;
  assign n1432 = n442 | n1431 ;
  assign n1433 = n290 & n1432 ;
  assign n1434 = n1430 | n1433 ;
  assign n1435 = n1420 & n1434 ;
  assign n1436 = n1406 | n1435 ;
  assign n1437 = ~n621 & n625 ;
  assign n1438 = ~n621 & n624 ;
  assign n1439 = n623 | n1438 ;
  assign n1440 = ~n1437 & n1439 ;
  assign n1441 = ~n75 & n1440 ;
  assign n1442 = ioin228 & n284 ;
  assign n1443 = ioin128 | n1442 ;
  assign n1444 = ioin228 & ioin128 ;
  assign n1445 = n291 & n1444 ;
  assign n1446 = n1443 & ~n1445 ;
  assign n1447 = n287 | n1446 ;
  assign n1448 = n287 & ~n1444 ;
  assign n1449 = n290 | n1448 ;
  assign n1450 = n1447 & ~n1449 ;
  assign n1451 = n283 | n1450 ;
  assign n1452 = n290 & n1418 ;
  assign n1453 = n1451 | n1452 ;
  assign n1454 = n283 & ~n1432 ;
  assign n1455 = n441 & ~n1454 ;
  assign n1456 = n1453 & n1455 ;
  assign n1457 = n1441 | n1456 ;
  assign n1458 = ~n617 & n619 ;
  assign n1459 = n582 & ~n1458 ;
  assign n1460 = ~n618 & n619 ;
  assign n1461 = n1459 | n1460 ;
  assign n1462 = ~n75 & n1461 ;
  assign n1463 = n283 & ~n1285 ;
  assign n1464 = n441 & ~n1463 ;
  assign n1465 = ioin227 & ioin127 ;
  assign n1466 = n287 & ~n1465 ;
  assign n1467 = n290 | n1466 ;
  assign n1468 = ioin227 & n284 ;
  assign n1469 = ioin127 | n1468 ;
  assign n1470 = n291 & n1465 ;
  assign n1471 = n1469 & ~n1470 ;
  assign n1472 = n287 | n1471 ;
  assign n1473 = ~n1467 & n1472 ;
  assign n1474 = n283 | n1473 ;
  assign n1475 = n290 & n1299 ;
  assign n1476 = n1474 | n1475 ;
  assign n1477 = n1464 & n1476 ;
  assign n1478 = n1462 | n1477 ;
  assign n1479 = n182 & ~n188 ;
  assign n1480 = n182 & ~n187 ;
  assign n1481 = n186 & ~n1480 ;
  assign n1482 = n1479 | n1481 ;
  assign n1483 = ~n75 & n1002 ;
  assign n1484 = n283 & ~n1190 ;
  assign n1485 = n441 & ~n1484 ;
  assign n1486 = ioin15 | n284 ;
  assign n1487 = ~n290 & n1486 ;
  assign n1488 = ioin15 & ~n287 ;
  assign n1489 = ioin25 & ~n1488 ;
  assign n1490 = ioin25 & n291 ;
  assign n1491 = n1488 & ~n1490 ;
  assign n1492 = n1489 | n1491 ;
  assign n1493 = n1487 & n1492 ;
  assign n1494 = n283 | n1493 ;
  assign n1495 = n290 & n1194 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n1485 & n1496 ;
  assign n1498 = n1483 | n1497 ;
  assign n1499 = ~n75 & n1055 ;
  assign n1500 = n283 & ~n437 ;
  assign n1501 = n441 & ~n1500 ;
  assign n1502 = ioin19 | n284 ;
  assign n1503 = ioin19 & ~n287 ;
  assign n1504 = ioin29 & ~n1503 ;
  assign n1505 = n1502 & n1504 ;
  assign n1506 = ioin29 & n291 ;
  assign n1507 = n1503 & ~n1506 ;
  assign n1508 = n1505 | n1507 ;
  assign n1509 = ~n290 & n1508 ;
  assign n1510 = n283 | n1509 ;
  assign n1511 = n290 & n476 ;
  assign n1512 = n1510 | n1511 ;
  assign n1513 = n1501 & n1512 ;
  assign n1514 = n1499 | n1513 ;
  assign n1515 = ~n75 & n1401 ;
  assign n1516 = n283 & ~n1153 ;
  assign n1517 = n441 & ~n1516 ;
  assign n1518 = ioin229 & n284 ;
  assign n1519 = ioin129 | n1518 ;
  assign n1520 = ioin229 & ioin129 ;
  assign n1521 = n291 & n1520 ;
  assign n1522 = n1519 & ~n1521 ;
  assign n1523 = n287 | n1522 ;
  assign n1524 = n287 & ~n1520 ;
  assign n1525 = n290 | n1524 ;
  assign n1526 = n1523 & ~n1525 ;
  assign n1527 = n283 | n1526 ;
  assign n1528 = n290 & n1167 ;
  assign n1529 = n1527 | n1528 ;
  assign n1530 = n1517 & n1529 ;
  assign n1531 = n1515 | n1530 ;
  assign n1532 = ~n75 & n1120 ;
  assign n1533 = ioin216 & ioin116 ;
  assign n1534 = n287 & ~n1533 ;
  assign n1535 = n290 | n1534 ;
  assign n1536 = ioin216 & n284 ;
  assign n1537 = ioin116 | n1536 ;
  assign n1538 = n291 & n1533 ;
  assign n1539 = n1537 & ~n1538 ;
  assign n1540 = n287 | n1539 ;
  assign n1541 = ~n1535 & n1540 ;
  assign n1542 = n283 | n1541 ;
  assign n1543 = n290 & n742 ;
  assign n1544 = n1542 | n1543 ;
  assign n1545 = n283 & ~n776 ;
  assign n1546 = n441 & ~n1545 ;
  assign n1547 = n1544 & n1546 ;
  assign n1548 = n1532 | n1547 ;
  assign n1549 = ~n75 & n1482 ;
  assign n1550 = n283 & ~n1379 ;
  assign n1551 = n441 & ~n1550 ;
  assign n1552 = ioin111 & ~n287 ;
  assign n1553 = ioin111 | n284 ;
  assign n1554 = ioin211 & n1553 ;
  assign n1555 = n1552 | n1554 ;
  assign n1556 = ioin211 & n291 ;
  assign n1557 = n1552 & n1556 ;
  assign n1558 = n290 | n1557 ;
  assign n1559 = n1555 & ~n1558 ;
  assign n1560 = n283 | n1559 ;
  assign n1561 = n290 & n1393 ;
  assign n1562 = n1560 | n1561 ;
  assign n1563 = n1551 & n1562 ;
  assign n1564 = n1549 | n1563 ;
  assign n1565 = ~n75 & n1219 ;
  assign n1566 = ioin16 & ioin26 ;
  assign n1567 = n287 & ~n1566 ;
  assign n1568 = n290 | n1567 ;
  assign n1569 = ioin26 & n284 ;
  assign n1570 = ioin16 | n1569 ;
  assign n1571 = n291 & n1566 ;
  assign n1572 = n1570 & ~n1571 ;
  assign n1573 = n287 | n1572 ;
  assign n1574 = ~n1568 & n1573 ;
  assign n1575 = n283 | n1574 ;
  assign n1576 = n290 & n865 ;
  assign n1577 = n1575 | n1576 ;
  assign n1578 = n283 & ~n901 ;
  assign n1579 = n441 & ~n1578 ;
  assign n1580 = n1577 & n1579 ;
  assign n1581 = n1565 | n1580 ;
  assign ioout22 = n480 ;
  assign ioadderout22 = n275 ;
  assign ioout7 = n560 ;
  assign iotestadderCout = n641 ;
  assign ioadderout17 = n645 ;
  assign ioadderout26 = n649 ;
  assign ioadderout1 = n653 ;
  assign ioadderout23 = n657 ;
  assign ioout1 = n723 ;
  assign ioadderout8 = n727 ;
  assign ioadderout0 = n729 ;
  assign ioadderout7 = n484 ;
  assign ioout15 = n780 ;
  assign ioout31 = n854 ;
  assign ioadderout10 = n858 ;
  assign ioout25 = n905 ;
  assign ioout10 = n948 ;
  assign ioout14 = n977 ;
  assign ioout24 = n998 ;
  assign ioadderout5 = n1002 ;
  assign ioout12 = n1051 ;
  assign ioadderout9 = n1055 ;
  assign ioadderout30 = n1059 ;
  assign ioadderout12 = n1006 ;
  assign ioadderout13 = n1063 ;
  assign ioout13 = n1095 ;
  assign ioout21 = n1116 ;
  assign ioadderout16 = n1120 ;
  assign ioout30 = n1136 ;
  assign ioadderout2 = n1140 ;
  assign ioout2 = n1171 ;
  assign ioadderout31 = n784 ;
  assign ioadderout14 = n952 ;
  assign ioout26 = n1198 ;
  assign ioout17 = n1215 ;
  assign ioadderout6 = n1219 ;
  assign ioout18 = n1240 ;
  assign ioout0 = n1266 ;
  assign ioout4 = n1303 ;
  assign ioout19 = n1324 ;
  assign ioadderout19 = n1307 ;
  assign ioout23 = n1349 ;
  assign ioout8 = n1365 ;
  assign ioadderout20 = n1369 ;
  assign ioout20 = n1397 ;
  assign ioadderout25 = n862 ;
  assign ioadderout29 = n1401 ;
  assign ioadderout15 = n733 ;
  assign ioout3 = n1436 ;
  assign ioout28 = n1457 ;
  assign ioout27 = n1478 ;
  assign ioadderout11 = n1482 ;
  assign ioout5 = n1498 ;
  assign ioadderout4 = n1270 ;
  assign ioout9 = n1514 ;
  assign ioadderout28 = n1440 ;
  assign ioadderout21 = n1114 ;
  assign ioadderout24 = n981 ;
  assign ioout29 = n1531 ;
  assign ioadderout27 = n1461 ;
  assign ioout16 = n1548 ;
  assign ioout11 = n1564 ;
  assign ioout6 = n1581 ;
  assign ioadderout3 = n1405 ;
  assign ioadderout18 = n1223 ;
endmodule
